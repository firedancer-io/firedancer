logic [385-1:0] out_p;
logic [385-1:0] out_n;
logic [M-1:0] p_m_o;
logic [M-1:0] n_m_o;
logic [4-1:0][M-1:0] p_m_o_p;
logic [415-1:0] p_s_1_00;
logic [294-1:0] p_s_0_00;
logic [287-1:0] p_s_0_06;
logic [265-1:0] p_s_0_18;
logic [294-1:0] p_s_0_12;
`SHADD_6_2C(294, p_s_0_00,   0,  10,  12,  24,  31,  33, {294'b0, in0[0+:260]}, {294'b0, in0[0+:260]}, {294'b0, in0[0+:260]}, {294'b0, in0[0+:260]}, {294'b0, in0[0+:260]}, {294'b0, in0[0+:260]});
`SHADD_6_2C(287, p_s_0_06,   0,   5,  10,  12,  15,  26, {287'b0, in0[0+:260]}, {287'b0, in0[0+:260]}, {287'b0, in0[0+:260]}, {287'b0, in0[0+:260]}, {287'b0, in0[0+:260]}, {287'b0, in0[0+:260]});
`SHADD_6_2C(294, p_s_0_12,   0,   5,  18,  21,  23,  33, {294'b0, in0[0+:260]}, {294'b0, in0[0+:260]}, {294'b0, in0[0+:260]}, {294'b0, in0[0+:260]}, {294'b0, in0[0+:260]}, {294'b0, in0[0+:260]});
`SHADD_6_2C(265, p_s_0_18,   0,   2,   4,   0,   0,   0, {265'b0, in0[0+:260]}, {265'b0, in0[0+:260]}, {265'b0, in0[0+:260]}, {265'b0, '0}, {265'b0, '0}, {265'b0, '0});
`SHADD_6_2C(415, p_s_1_00,   0,  37,  72, 120,   0,   0, {415'b0, p_s_0_00}, {415'b0, p_s_0_06}, {415'b0, p_s_0_12}, {415'b0, p_s_0_18}, {415'b0, '0}, {415'b0, '0});
assign out_p = p_s_1_00 << 0;
assign p_m_o = p_m_o_p[4-1];
always_ff@(posedge clk) p_m_o_p[0] <= m_i;
always_ff@(posedge clk) p_m_o_p[1] <= p_m_o_p[1-1];
always_ff@(posedge clk) p_m_o_p[2] <= p_m_o_p[2-1];
always_ff@(posedge clk) p_m_o_p[3] <= p_m_o_p[3-1];
logic [4-1:0][M-1:0] n_m_o_p;
logic [293-1:0] n_s_0_06;
logic [380-1:0] n_s_1_00;
logic [285-1:0] n_s_0_00;
logic [279-1:0] n_s_0_12;
logic [290-1:0] n_s_0_18;
`SHADD_6_2C(285, n_s_0_00,   0,   2,  12,  15,  17,  24, {285'b0, in0[0+:260]}, {285'b0, in0[0+:260]}, {285'b0, in0[0+:260]}, {285'b0, in0[0+:260]}, {285'b0, in0[0+:260]}, {285'b0, in0[0+:260]});
`SHADD_6_2C(293, n_s_0_06,   0,   6,  11,  16,  30,  32, {293'b0, in0[0+:260]}, {293'b0, in0[0+:260]}, {293'b0, in0[0+:260]}, {293'b0, in0[0+:260]}, {293'b0, in0[0+:260]}, {293'b0, in0[0+:260]});
`SHADD_6_2C(279, n_s_0_12,   0,   2,   4,   9,  14,  18, {279'b0, in0[0+:260]}, {279'b0, in0[0+:260]}, {279'b0, in0[0+:260]}, {279'b0, in0[0+:260]}, {279'b0, in0[0+:260]}, {279'b0, in0[0+:260]});
`SHADD_6_2C(290, n_s_0_18,   0,   9,  13,  19,  24,  29, {290'b0, in0[0+:260]}, {290'b0, in0[0+:260]}, {290'b0, in0[0+:260]}, {290'b0, in0[0+:260]}, {290'b0, in0[0+:260]}, {290'b0, in0[0+:260]});
`SHADD_6_2C(380, n_s_1_00,   0,  27,  63,  86,   0,   0, {380'b0, n_s_0_00}, {380'b0, n_s_0_06}, {380'b0, n_s_0_12}, {380'b0, n_s_0_18}, {380'b0, '0}, {380'b0, '0});
assign out_n = n_s_1_00 << 2;
assign n_m_o = n_m_o_p[4-1];
always_ff@(posedge clk) n_m_o_p[0] <= m_i;
always_ff@(posedge clk) n_m_o_p[1] <= n_m_o_p[1-1];
always_ff@(posedge clk) n_m_o_p[2] <= n_m_o_p[2-1];
always_ff@(posedge clk) n_m_o_p[3] <= n_m_o_p[3-1];
always_ff@(posedge clk) out0 <= out_p - out_n;
always_ff@(posedge clk) m_o <= p_m_o;
